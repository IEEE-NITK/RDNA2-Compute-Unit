`include "VOP2.sv"
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: IEEE NITK
// Engineer: Kruti Deepan Panda
// 
// Create Date: 04.10.2021 18:48:26
// Design Name: ALU
// Module Name: VOP2_ALU
// Project Name: RDNA2 Compute Unit 
//////////////////////////////////////////////////////////////////////////////////


module VOP2_ALU(
input wire instruction[31:0]
    );
    
endmodule
