`ifndef _scalars_vh
`define _scalars_vh

//Scalar instruction constants
localparam SOP1 = 7'b1111101;
localparam SOPK = 2'b11;
localparam SOPC=7'b1111110

`endif