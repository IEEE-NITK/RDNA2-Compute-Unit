`ifndef _trial_vh
`define _trial_vh

//32 bit constants for floating point numbers
localparam pos_inf_32 = 32'b01111111100000000000000000000000;

`endif
