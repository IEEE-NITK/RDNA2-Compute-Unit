`ifndef VOP2
`define VOP2

`define V_ADD_F16       	 	32'b0
`define V_ADD_F32       	 	32'b0
`define V_ADD_CO_CI_U32			32'b0
`define V_ADD_NC_U32			32'b0
`define V_AND_B32    			32'b0
`define V_ASHRREV_B32			32'b0
`define V_CNDMASK_B32 			32'b0
`define V_CVT_PKRTZ_F16_F32		32'b0
`define V_FMAAK_F16 			32'b0
`define V_FMAAK_F32			    32'b0
`define V_FMAC_F16			    32'b0
`define V_FMAC_F32			    32'b0
`define V_FMAMK_F16			    32'b0
`define V_FMAMK_F32 			32'b0
`define V_LDEXP_F16 			32'b0
`define V_LSHLREV_B32			32'b0
`define V_LSHRREV_B32 			32'b0
`define V_MAC_{ F16,F32} 		32'b0
`define V_MAX_{ F16, F32,I32,U32} 	32'b0
`define V_MIN_{ F16, F32,I32,U32} 	32'b0
`define V_MUL_F16       		32'b0
`define V_MUL_F32       		32'b0
`define V_MUL_HI_I32_I24		32'b0
`define V_MUL_HI_U32_U24		32'b0
`define V_MUL_I32_I24 			32'b0
`define V_MUL_LEGACY_F32		32'b0
`define V_MUL_U32_U24			32'b0
`define V_OR_B32		      	32'b0
`define V_SUB_F16        		32'b0
`define V_SUB_F32        		32'b0
`define V_SUB_CO_CI_U32			32'b0
`define V_SUB_NC_U32			32'b0
`define V_SUBREV_F16    		32'b0
`define V_SUBREV_F32    		32'b0
`define V_SUBREV_CO_CI_U32		32'b0
`define V_SUBREV_NC_U32			32'b0
`define V_XNOR_B32  			32'b0
`define V_XOR_B32    			32'b0
`define V_DOT2C_F32_F16 		32'b0
`define V_DOT4C_I32_I8			32'b0

`endif
