`ifndef _scalars_vh
`define _scalars_vh

//Scalar instruction constants
localparam SOP1 = 7'b1111101;


`endif