`include "floats.vh"
`timescale 1ns / 1ps


module float_adder_32(
    input [31:0] A,
    input [31:0] B,
    output [31:0] out
    );
endmodule
